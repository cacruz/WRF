netcdf force_template {
dimensions:
	Time = UNLIMITED ; // (0 currently)
	DateStrLen = 19 ;
	force_layers = 29 ;
variables:
	char Times(Time, DateStrLen) ;
	float Z_FORCE(Time, force_layers) ;
		Z_FORCE:FieldType = 104 ;
		Z_FORCE:MemoryOrder = "Z  " ;
		Z_FORCE:description = "height of forcing time series" ;
		Z_FORCE:units = "" ;
		Z_FORCE:stagger = "" ;
		Z_FORCE:_FillValue = -999.f ;
	float Z_FORCE_TEND(Time, force_layers) ;
		Z_FORCE_TEND:FieldType = 104 ;
		Z_FORCE_TEND:MemoryOrder = "Z  " ;
		Z_FORCE_TEND:description = "tendency height of forcing time series" ;
		Z_FORCE_TEND:units = "" ;
		Z_FORCE_TEND:stagger = "" ;
		Z_FORCE_TEND:_FillValue = -999.f ;
	float U_G(Time, force_layers) ;
		U_G:FieldType = 104 ;
		U_G:MemoryOrder = "Z  " ;
		U_G:description = "x-component geostrophic wind" ;
		U_G:units = "m s-1" ;
		U_G:stagger = "" ;
		U_G:_FillValue = -999.f ;
	float U_G_TEND(Time, force_layers) ;
		U_G_TEND:FieldType = 104 ;
		U_G_TEND:MemoryOrder = "Z  " ;
		U_G_TEND:description = "tendency x-component geostrophic wind" ;
		U_G_TEND:units = "m s-2" ;
		U_G_TEND:stagger = "" ;
	float V_G(Time, force_layers) ;
		V_G:FieldType = 104 ;
		V_G:MemoryOrder = "Z  " ;
		V_G:description = "y-component geostrophic wind" ;
		V_G:units = "m s-1" ;
		V_G:stagger = "" ;
		V_G:_FillValue = -999.f ;
	float V_G_TEND(Time, force_layers) ;
		V_G_TEND:FieldType = 104 ;
		V_G_TEND:MemoryOrder = "Z  " ;
		V_G_TEND:description = "tendency y-component geostrophic wind" ;
		V_G_TEND:units = "m s-2" ;
		V_G_TEND:stagger = "" ;
	float W_SUBS(Time, force_layers) ;
		W_SUBS:FieldType = 104 ;
		W_SUBS:MemoryOrder = "Z  " ;
		W_SUBS:description = "large-scale vertical motion (subsidence)" ;
		W_SUBS:units = "m s-1" ;
		W_SUBS:stagger = "" ;
		W_SUBS:_FillValue = -999.f ;
	float W_SUBS_TEND(Time, force_layers) ;
		W_SUBS_TEND:FieldType = 104 ;
		W_SUBS_TEND:MemoryOrder = "Z  " ;
		W_SUBS_TEND:description = "tendency large-scale vertical motion (subsidence)" ;
		W_SUBS_TEND:units = "m s-2" ;
		W_SUBS_TEND:stagger = "" ;
	float TH_UPSTREAM_X(Time, force_layers) ;
		TH_UPSTREAM_X:FieldType = 104 ;
		TH_UPSTREAM_X:MemoryOrder = "Z  " ;
		TH_UPSTREAM_X:description = "upstream theta x-advection" ;
		TH_UPSTREAM_X:units = "K s-1" ;
		TH_UPSTREAM_X:stagger = "" ;
	float TH_UPSTREAM_X_TEND(Time, force_layers) ;
		TH_UPSTREAM_X_TEND:FieldType = 104 ;
		TH_UPSTREAM_X_TEND:MemoryOrder = "Z  " ;
		TH_UPSTREAM_X_TEND:description = "tendency upstream theta x-advection" ;
		TH_UPSTREAM_X_TEND:units = "K s-2" ;
		TH_UPSTREAM_X_TEND:stagger = "" ;
	float TH_UPSTREAM_Y(Time, force_layers) ;
		TH_UPSTREAM_Y:FieldType = 104 ;
		TH_UPSTREAM_Y:MemoryOrder = "Z  " ;
		TH_UPSTREAM_Y:description = "upstream theta y-advection" ;
		TH_UPSTREAM_Y:units = "K s-1" ;
		TH_UPSTREAM_Y:stagger = "" ;
	float TH_UPSTREAM_Y_TEND(Time, force_layers) ;
		TH_UPSTREAM_Y_TEND:FieldType = 104 ;
		TH_UPSTREAM_Y_TEND:MemoryOrder = "Z  " ;
		TH_UPSTREAM_Y_TEND:description = "tendency upstream theta y-advection" ;
		TH_UPSTREAM_Y_TEND:units = "K s-2" ;
		TH_UPSTREAM_Y_TEND:stagger = "" ;
	float QV_UPSTREAM_X(Time, force_layers) ;
		QV_UPSTREAM_X:FieldType = 104 ;
		QV_UPSTREAM_X:MemoryOrder = "Z  " ;
		QV_UPSTREAM_X:description = "upstream qv x-advection" ;
		QV_UPSTREAM_X:units = "kg kg-1 s-1" ;
		QV_UPSTREAM_X:stagger = "" ;
	float QV_UPSTREAM_X_TEND(Time, force_layers) ;
		QV_UPSTREAM_X_TEND:FieldType = 104 ;
		QV_UPSTREAM_X_TEND:MemoryOrder = "Z  " ;
		QV_UPSTREAM_X_TEND:description = "tendency upstream qv x-advection" ;
		QV_UPSTREAM_X_TEND:units = "kg kg-1 s-2" ;
		QV_UPSTREAM_X_TEND:stagger = "" ;
	float QV_UPSTREAM_Y(Time, force_layers) ;
		QV_UPSTREAM_Y:FieldType = 104 ;
		QV_UPSTREAM_Y:MemoryOrder = "Z  " ;
		QV_UPSTREAM_Y:description = "upstream qv y-advection" ;
		QV_UPSTREAM_Y:units = "kg kg-1 s-1" ;
		QV_UPSTREAM_Y:stagger = "" ;
	float QV_UPSTREAM_Y_TEND(Time, force_layers) ;
		QV_UPSTREAM_Y_TEND:FieldType = 104 ;
		QV_UPSTREAM_Y_TEND:MemoryOrder = "Z  " ;
		QV_UPSTREAM_Y_TEND:description = "tendency upstream qv y-advection" ;
		QV_UPSTREAM_Y_TEND:units = "kg kg-1 s-2" ;
		QV_UPSTREAM_Y_TEND:stagger = "" ;
	float U_UPSTREAM_X(Time, force_layers) ;
		U_UPSTREAM_X:FieldType = 104 ;
		U_UPSTREAM_X:MemoryOrder = "Z  " ;
		U_UPSTREAM_X:description = "upstream U x-advection" ;
		U_UPSTREAM_X:units = "m s-3" ;
		U_UPSTREAM_X:stagger = "" ;
	float U_UPSTREAM_X_TEND(Time, force_layers) ;
		U_UPSTREAM_X_TEND:FieldType = 104 ;
		U_UPSTREAM_X_TEND:MemoryOrder = "Z  " ;
		U_UPSTREAM_X_TEND:description = "tendency upstream U x-advection" ;
		U_UPSTREAM_X_TEND:units = "m s-3" ;
		U_UPSTREAM_X_TEND:stagger = "" ;
	float U_UPSTREAM_Y(Time, force_layers) ;
		U_UPSTREAM_Y:FieldType = 104 ;
		U_UPSTREAM_Y:MemoryOrder = "Z  " ;
		U_UPSTREAM_Y:description = "upstream U y-advection" ;
		U_UPSTREAM_Y:units = "m s-3" ;
		U_UPSTREAM_Y:stagger = "" ;
	float U_UPSTREAM_Y_TEND(Time, force_layers) ;
		U_UPSTREAM_Y_TEND:FieldType = 104 ;
		U_UPSTREAM_Y_TEND:MemoryOrder = "Z  " ;
		U_UPSTREAM_Y_TEND:description = "tendency upstream U y-advection" ;
		U_UPSTREAM_Y_TEND:units = "m s-3" ;
		U_UPSTREAM_Y_TEND:stagger = "" ;
	float V_UPSTREAM_X(Time, force_layers) ;
		V_UPSTREAM_X:FieldType = 104 ;
		V_UPSTREAM_X:MemoryOrder = "Z  " ;
		V_UPSTREAM_X:description = "upstream V x-advection" ;
		V_UPSTREAM_X:units = "m s-3" ;
		V_UPSTREAM_X:stagger = "" ;
	float V_UPSTREAM_X_TEND(Time, force_layers) ;
		V_UPSTREAM_X_TEND:FieldType = 104 ;
		V_UPSTREAM_X_TEND:MemoryOrder = "Z  " ;
		V_UPSTREAM_X_TEND:description = "tendency upstream V x-advection" ;
		V_UPSTREAM_X_TEND:units = "m s-3" ;
		V_UPSTREAM_X_TEND:stagger = "" ;
	float V_UPSTREAM_Y(Time, force_layers) ;
		V_UPSTREAM_Y:FieldType = 104 ;
		V_UPSTREAM_Y:MemoryOrder = "Z  " ;
		V_UPSTREAM_Y:description = "upstream V y-advection" ;
		V_UPSTREAM_Y:units = "m s-3" ;
		V_UPSTREAM_Y:stagger = "" ;
	float V_UPSTREAM_Y_TEND(Time, force_layers) ;
		V_UPSTREAM_Y_TEND:FieldType = 104 ;
		V_UPSTREAM_Y_TEND:MemoryOrder = "Z  " ;
		V_UPSTREAM_Y_TEND:description = "tendency upstream V y-advection" ;
		V_UPSTREAM_Y_TEND:units = "m s-3" ;
		V_UPSTREAM_Y_TEND:stagger = "" ;
	float TAU_X(Time, force_layers) ;
		TAU_X:FieldType = 104 ;
		TAU_X:MemoryOrder = "Z  " ;
		TAU_X:description = "X-direction advective timescale" ;
		TAU_X:units = "s" ;
		TAU_X:stagger = "" ;
	float TAU_X_TEND(Time, force_layers) ;
		TAU_X_TEND:FieldType = 104 ;
		TAU_X_TEND:MemoryOrder = "Z  " ;
		TAU_X_TEND:description = "tendency X-direction advective timescale" ;
		TAU_X_TEND:units = "" ;
		TAU_X_TEND:stagger = "" ;
	float TAU_Y(Time, force_layers) ;
		TAU_Y:FieldType = 104 ;
		TAU_Y:MemoryOrder = "Z  " ;
		TAU_Y:description = "Y-direction advective timescale" ;
		TAU_Y:units = "s" ;
		TAU_Y:stagger = "" ;
	float TAU_Y_TEND(Time, force_layers) ;
		TAU_Y_TEND:FieldType = 104 ;
		TAU_Y_TEND:MemoryOrder = "Z  " ;
		TAU_Y_TEND:description = "tendency Y-direction advective timescale" ;
		TAU_Y_TEND:units = "" ;
		TAU_Y_TEND:stagger = "" ;

// global attributes:
		:TITLE = "AUXILIARY FORCING FOR SCM" ;
		:START_DATE = "2003-05-03_12:00:00" ;
		:SIMULATION_START_DATE = "2003-05-03_12:00:00" ;
		:DX = 4000.f ;
		:DY = 4000.f ;
		:GRID_ID = 1 ;
		:PARENT_ID = 0 ;
		:I_PARENT_START = 1 ;
		:J_PARENT_START = 1 ;
		:PARENT_GRID_RATIO = 1 ;
		:DT = 20.f ;
		:CEN_LAT = 0.f ;
		:CEN_LON = 0.f ;
		:TRUELAT1 = 0.f ;
		:TRUELAT2 = 0.f ;
		:MOAD_CEN_LAT = 0.f ;
		:STAND_LON = 0.f ;
		:GMT = 0.f ;
		:JULYR = 0 ;
		:JULDAY = 1 ;
		:MAP_PROJ = 0 ;
		:MMINLU = "USGS" ;
		:ISWATER = 16 ;
		:ISICE = 0 ;
		:ISURBAN = 0 ;
		:ISOILWATER = 0 ;
}
